module extend (
	Instr,
	ImmSrc,
	ExtImm
);
	input wire [23:0] Instr;
	input wire [1:0] ImmSrc;
	output reg [31:0] ExtImm;
	always @(*)
		case (ImmSrc)
			2'b00: ExtImm = {24'b000000000000000000000000, Instr[7:0]}; // Imm8
			2'b01: ExtImm = {20'b00000000000000000000, Instr[11:0]}; // Imm12
			2'b10: ExtImm = {{6 {Instr[23]}}, Instr[23:0], 2'b00}; // Imm24 (con bit extension)
			default: ExtImm = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
		endcase
endmodule